module top (
    input         clk,
    input         n_rst,
    input   [7:0] data_in,
    output  [7:0] data_out,
    input  [15:0] address_out
);

endmodule
