module cpu (
    input clk, 
    input reset
);

endmodule;
